// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 18.0.0 Build 614 04/24/2018 SJ Lite Edition"
// CREATED		"Tue May 29 15:02:09 2018"

module serializer(
	CLOCK_50,
	serial
);


input wire	CLOCK_50;
output wire	serial;

wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	[7:0] SYNTHESIZED_WIRE_3;





baud_clock	b2v_inst(
	.inclk0(CLOCK_50),
	.c0(SYNTHESIZED_WIRE_6));


down_count	b2v_inst1(
	.clock(SYNTHESIZED_WIRE_5),
	.q(SYNTHESIZED_WIRE_3));


serialize	b2v_inst3(
	.send(SYNTHESIZED_WIRE_5),
	.baud(SYNTHESIZED_WIRE_6),
	.count(SYNTHESIZED_WIRE_3),
	.out(serial));


send_data	b2v_inst5(
	.clk(SYNTHESIZED_WIRE_6),
	.tick(SYNTHESIZED_WIRE_5));


endmodule
